* SPICE3 file created from inv_std_layout.ext - technology: scmos

M1000 Out in Gnd Gnd nfet w=1.2u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
M1001 Out in Vdd Vdd pfet w=2u l=0.4u
+  ad=0p pd=0u as=0p ps=0u
C0 Out in 0.04fF
C1 Vdd Out 0.23fF
C2 Vdd in 0.34fF
C3 Out Gnd 0.10fF
C4 in Gnd 0.23fF
C5 Vdd Gnd 1.66fF

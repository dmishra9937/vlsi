magic
tech scmos
timestamp 1661171676
<< nwell >>
rect -16 -2 31 19
<< ntransistor >>
rect 6 -18 9 -11
<< ptransistor >>
rect 6 5 9 13
<< ndiffusion >>
rect 2 -18 6 -11
rect 9 -18 17 -11
<< pdiffusion >>
rect 1 5 6 13
rect 9 5 17 13
<< ndcontact >>
rect -2 -18 2 -11
rect 17 -18 21 -11
<< pdcontact >>
rect -3 5 1 13
rect 17 5 21 13
<< psubstratepcontact >>
rect -10 -18 -6 -11
<< nsubstratencontact >>
rect -11 5 -7 13
<< polysilicon >>
rect 6 13 9 15
rect 6 2 9 5
rect 8 -2 9 2
rect 6 -11 9 -2
rect 6 -20 9 -18
<< polycontact >>
rect 4 -2 8 2
<< metal1 >>
rect -11 16 20 19
rect -7 5 -3 16
rect 1 -2 4 1
rect 8 -2 9 1
rect 18 -11 21 5
rect -6 -25 -2 -11
rect -9 -28 22 -25
<< labels >>
rlabel metal1 -6 17 -6 17 5 vdd
rlabel metal1 -5 -26 -5 -26 1 gnd
rlabel metal1 3 0 3 0 1 in
rlabel metal1 19 -4 19 -4 1 out
<< end >>

magic
tech scmos
timestamp 1661604029
<< nwell >>
rect -3 3 32 25
<< ntransistor >>
rect 9 -9 11 -3
rect 17 -9 19 -3
<< ptransistor >>
rect 9 9 11 19
rect 17 9 19 19
<< ndiffusion >>
rect 1 -4 9 -3
rect 1 -8 4 -4
rect 8 -8 9 -4
rect 1 -9 9 -8
rect 11 -4 17 -3
rect 11 -8 12 -4
rect 16 -8 17 -4
rect 11 -9 17 -8
rect 19 -4 27 -3
rect 19 -8 21 -4
rect 25 -8 27 -4
rect 19 -9 27 -8
<< pdiffusion >>
rect 3 18 9 19
rect 3 10 4 18
rect 8 10 9 18
rect 3 9 9 10
rect 11 18 17 19
rect 11 10 12 18
rect 16 10 17 18
rect 11 9 17 10
rect 19 18 25 19
rect 19 10 20 18
rect 24 10 25 18
rect 19 9 25 10
<< ndcontact >>
rect 4 -8 8 -4
rect 12 -8 16 -4
rect 21 -8 25 -4
<< pdcontact >>
rect 4 10 8 18
rect 12 10 16 18
rect 20 10 24 18
<< polysilicon >>
rect 9 19 11 21
rect 17 19 19 21
rect 9 5 11 9
rect 9 -3 11 1
rect 17 -3 19 9
rect 9 -11 11 -9
rect 17 -11 19 -9
<< polycontact >>
rect 6 1 11 5
<< metal1 >>
rect 3 22 11 25
rect 4 18 8 22
rect 4 9 8 10
rect 3 1 6 5
rect 4 -4 8 -3
rect 21 -4 25 -3
rect 4 -12 8 -8
rect 21 -12 25 -8
rect 2 -15 26 -12
<< metal2 >>
rect 20 5 24 19
rect 12 2 28 5
rect 12 -9 16 2
<< labels >>
rlabel metal1 6 23 6 23 5 Vdd!
rlabel metal2 25 3 25 3 1 Out
rlabel metal1 13 -14 13 -14 1 gnd!
rlabel metal1 5 3 5 3 1 In
<< end >>
